Library ieee;
Use ieee.std_logic_1164.all;

entity ExecuteStage is
  port (
    clock:IN std_logic
  ) ;
end ExecuteStage;