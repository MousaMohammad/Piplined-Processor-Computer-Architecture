Library ieee;
Use ieee.std_logic_1164.all;

entity ExMem_buf is
  port (
    Rst, Clk : IN STD_LOGIC;
    -- Ex ports --
    
  );
end entity;

architecture arch of ExMem_buf is
begin

end arch ; -- arch
