Library ieee;
Use ieee.std_logic_1164.all;

entity ExWB_buf is
  port (
    Rst, Clk : IN STD_LOGIC
  ) ;
end ExWB_buf;


architecture archbuf of ExWB_buf is 

begin

end archbuf ; -- archbuf


